`include "am2940_interface.sv"
`include "am2940_base_unit.sv"
`include "am2940_packet.sv"
`include "am2940_data_in_generator.sv"
`include "am2940_data_in_bfm.sv"
`include "am2940_address_out_generator.sv"
`include "am2940_address_out_bfm.sv"
`include "am2940_data_in_monitor.sv"
`include "am2940_address_out_monitor.sv"
`include "am2940_sb.sv"
`include "am2940_environment.sv"